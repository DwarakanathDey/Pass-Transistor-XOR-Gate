module dwaraka_NOT (output Y, input A);
    not (Y, A);
endmodule
